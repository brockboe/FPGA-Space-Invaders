// sprite_rom.sv
//
// stores data about enemy sprites

module sprite_rom
(
	input 	[7:0] addr,
	output 	[7:0] data
);

	logic[7:0] addr_reg;

	parameter [0:48][7:0] ROM = {

		8'b01000010, //0  █    █ 
		8'b00100100, //1   █  █  
		8'b01011010, //2  █ ██ █ 
		8'b11111111, //3 ████████
		8'b10100101, //4 █ █  █ █
		8'b00011000, //5    ██   
		8'b00000000, //6 
		8'b00000000, //7 
		
		8'b00100100, //8    █  █  
		8'b00100100, //9    █  █  
		8'b01011010, //10  █ ██ █
		8'b11111111, //11 ████████
		8'b10100101, //12 █ █  █ █
		8'b00100100, //13   █  █  
		8'b01000010, //14  █    █
		8'b00000000, //15 
		
		8'b00011000, //16    ██   
		8'b00111100, //17   ████  
		8'b01111110, //18  ██████
		8'b01101010, //19  ██ █ █
		8'b01111110, //20  ██████
		8'b01111110, //21  ██████
		8'b00101010, //22   █ █ █
		8'b00000000, //23
		
		8'b00011000, //24    ██   
		8'b00111100, //25   ████  
		8'b01111110, //26  ██████ 
		8'b01010110, //27  █ █ ██
		8'b01111110, //28  ██████
		8'b01111110, //29  ██████
		8'b01010100, //30  █ █ █ 
		8'b00000000, //31
		
		8'b00111100, //32   ████  
		8'b01111110, //33  ██████ 
		8'b10011001, //34 █  ██  █
		8'b11111111, //35 ████████
		8'b00000000, //36 
		8'b01100110, //37  ██  ██
		8'b10011001, //38 █  ██  █
		8'b00000000, //39 
		
		8'b00111100, //40   ████  
		8'b01111110, //41  ██████ 
		8'b11011011, //42 ██ ██ ██
		8'b11111111, //43 ████████
		8'b00000000, //44
		8'b00100100, //45   █  █  
		8'b11011011, //46 ██ ██ ██
		8'b00000000  //47
		
	};

	assign data = ROM[addr];
	
endmodule 